client jjAIS
is
	interface jiAIS;
end ;