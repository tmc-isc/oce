interface jiAIS
is
	package AIS;
end ;